`timescale 1ns / 1ps

module Adder(SUM,A,B);
		input A,B;
		output SUM;
		assign SUM = A + B;
endmodule
